module top_module (
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);//

    add16 first (  );
    add16 secnd (  );
    
endmodule

module add1 ( input a, input b, input cin,   output sum, output cout );

// Full adder module here

endmodule